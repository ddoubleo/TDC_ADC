module TDC ( 
 input clk, 
 input start, 
 output [254:0] regs_out,
 output out
);

wire out0 /* synthesis syn_keep=1 */ ;
wire out1 /* synthesis syn_keep=1 */ ;
wire out2 /* synthesis syn_keep=1 */ ;
wire out3 /* synthesis syn_keep=1 */ ;
wire out4 /* synthesis syn_keep=1 */ ;
wire out5 /* synthesis syn_keep=1 */ ;
wire out6 /* synthesis syn_keep=1 */ ;
wire out7 /* synthesis syn_keep=1 */ ;
wire out8 /* synthesis syn_keep=1 */ ;
wire out9 /* synthesis syn_keep=1 */ ;
wire out10 /* synthesis syn_keep=1 */ ;
wire out11 /* synthesis syn_keep=1 */ ;
wire out12 /* synthesis syn_keep=1 */ ;
wire out13 /* synthesis syn_keep=1 */ ;
wire out14 /* synthesis syn_keep=1 */ ;
wire out15 /* synthesis syn_keep=1 */ ;
wire out16 /* synthesis syn_keep=1 */ ;
wire out17 /* synthesis syn_keep=1 */ ;
wire out18 /* synthesis syn_keep=1 */ ;
wire out19 /* synthesis syn_keep=1 */ ;
wire out20 /* synthesis syn_keep=1 */ ;
wire out21 /* synthesis syn_keep=1 */ ;
wire out22 /* synthesis syn_keep=1 */ ;
wire out23 /* synthesis syn_keep=1 */ ;
wire out24 /* synthesis syn_keep=1 */ ;
wire out25 /* synthesis syn_keep=1 */ ;
wire out26 /* synthesis syn_keep=1 */ ;
wire out27 /* synthesis syn_keep=1 */ ;
wire out28 /* synthesis syn_keep=1 */ ;
wire out29 /* synthesis syn_keep=1 */ ;
wire out30 /* synthesis syn_keep=1 */ ;
wire out31 /* synthesis syn_keep=1 */ ;
wire out32 /* synthesis syn_keep=1 */ ;
wire out33 /* synthesis syn_keep=1 */ ;
wire out34 /* synthesis syn_keep=1 */ ;
wire out35 /* synthesis syn_keep=1 */ ;
wire out36 /* synthesis syn_keep=1 */ ;
wire out37 /* synthesis syn_keep=1 */ ;
wire out38 /* synthesis syn_keep=1 */ ;
wire out39 /* synthesis syn_keep=1 */ ;
wire out40 /* synthesis syn_keep=1 */ ;
wire out41 /* synthesis syn_keep=1 */ ;
wire out42 /* synthesis syn_keep=1 */ ;
wire out43 /* synthesis syn_keep=1 */ ;
wire out44 /* synthesis syn_keep=1 */ ;
wire out45 /* synthesis syn_keep=1 */ ;
wire out46 /* synthesis syn_keep=1 */ ;
wire out47 /* synthesis syn_keep=1 */ ;
wire out48 /* synthesis syn_keep=1 */ ;
wire out49 /* synthesis syn_keep=1 */ ;
wire out50 /* synthesis syn_keep=1 */ ;
wire out51 /* synthesis syn_keep=1 */ ;
wire out52 /* synthesis syn_keep=1 */ ;
wire out53 /* synthesis syn_keep=1 */ ;
wire out54 /* synthesis syn_keep=1 */ ;
wire out55 /* synthesis syn_keep=1 */ ;
wire out56 /* synthesis syn_keep=1 */ ;
wire out57 /* synthesis syn_keep=1 */ ;
wire out58 /* synthesis syn_keep=1 */ ;
wire out59 /* synthesis syn_keep=1 */ ;
wire out60 /* synthesis syn_keep=1 */ ;
wire out61 /* synthesis syn_keep=1 */ ;
wire out62 /* synthesis syn_keep=1 */ ;
wire out63 /* synthesis syn_keep=1 */ ;
wire out64 /* synthesis syn_keep=1 */ ;
wire out65 /* synthesis syn_keep=1 */ ;
wire out66 /* synthesis syn_keep=1 */ ;
wire out67 /* synthesis syn_keep=1 */ ;
wire out68 /* synthesis syn_keep=1 */ ;
wire out69 /* synthesis syn_keep=1 */ ;
wire out70 /* synthesis syn_keep=1 */ ;
wire out71 /* synthesis syn_keep=1 */ ;
wire out72 /* synthesis syn_keep=1 */ ;
wire out73 /* synthesis syn_keep=1 */ ;
wire out74 /* synthesis syn_keep=1 */ ;
wire out75 /* synthesis syn_keep=1 */ ;
wire out76 /* synthesis syn_keep=1 */ ;
wire out77 /* synthesis syn_keep=1 */ ;
wire out78 /* synthesis syn_keep=1 */ ;
wire out79 /* synthesis syn_keep=1 */ ;
wire out80 /* synthesis syn_keep=1 */ ;
wire out81 /* synthesis syn_keep=1 */ ;
wire out82 /* synthesis syn_keep=1 */ ;
wire out83 /* synthesis syn_keep=1 */ ;
wire out84 /* synthesis syn_keep=1 */ ;
wire out85 /* synthesis syn_keep=1 */ ;
wire out86 /* synthesis syn_keep=1 */ ;
wire out87 /* synthesis syn_keep=1 */ ;
wire out88 /* synthesis syn_keep=1 */ ;
wire out89 /* synthesis syn_keep=1 */ ;
wire out90 /* synthesis syn_keep=1 */ ;
wire out91 /* synthesis syn_keep=1 */ ;
wire out92 /* synthesis syn_keep=1 */ ;
wire out93 /* synthesis syn_keep=1 */ ;
wire out94 /* synthesis syn_keep=1 */ ;
wire out95 /* synthesis syn_keep=1 */ ;
wire out96 /* synthesis syn_keep=1 */ ;
wire out97 /* synthesis syn_keep=1 */ ;
wire out98 /* synthesis syn_keep=1 */ ;
wire out99 /* synthesis syn_keep=1 */ ;
wire out100 /* synthesis syn_keep=1 */ ;
wire out101 /* synthesis syn_keep=1 */ ;
wire out102 /* synthesis syn_keep=1 */ ;
wire out103 /* synthesis syn_keep=1 */ ;
wire out104 /* synthesis syn_keep=1 */ ;
wire out105 /* synthesis syn_keep=1 */ ;
wire out106 /* synthesis syn_keep=1 */ ;
wire out107 /* synthesis syn_keep=1 */ ;
wire out108 /* synthesis syn_keep=1 */ ;
wire out109 /* synthesis syn_keep=1 */ ;
wire out110 /* synthesis syn_keep=1 */ ;
wire out111 /* synthesis syn_keep=1 */ ;
wire out112 /* synthesis syn_keep=1 */ ;
wire out113 /* synthesis syn_keep=1 */ ;
wire out114 /* synthesis syn_keep=1 */ ;
wire out115 /* synthesis syn_keep=1 */ ;
wire out116 /* synthesis syn_keep=1 */ ;
wire out117 /* synthesis syn_keep=1 */ ;
wire out118 /* synthesis syn_keep=1 */ ;
wire out119 /* synthesis syn_keep=1 */ ;
wire out120 /* synthesis syn_keep=1 */ ;
wire out121 /* synthesis syn_keep=1 */ ;
wire out122 /* synthesis syn_keep=1 */ ;
wire out123 /* synthesis syn_keep=1 */ ;
wire out124 /* synthesis syn_keep=1 */ ;
wire out125 /* synthesis syn_keep=1 */ ;
wire out126 /* synthesis syn_keep=1 */ ;
wire out127 /* synthesis syn_keep=1 */ ;
wire out128 /* synthesis syn_keep=1 */ ;
wire out129 /* synthesis syn_keep=1 */ ;
wire out130 /* synthesis syn_keep=1 */ ;
wire out131 /* synthesis syn_keep=1 */ ;
wire out132 /* synthesis syn_keep=1 */ ;
wire out133 /* synthesis syn_keep=1 */ ;
wire out134 /* synthesis syn_keep=1 */ ;
wire out135 /* synthesis syn_keep=1 */ ;
wire out136 /* synthesis syn_keep=1 */ ;
wire out137 /* synthesis syn_keep=1 */ ;
wire out138 /* synthesis syn_keep=1 */ ;
wire out139 /* synthesis syn_keep=1 */ ;
wire out140 /* synthesis syn_keep=1 */ ;
wire out141 /* synthesis syn_keep=1 */ ;
wire out142 /* synthesis syn_keep=1 */ ;
wire out143 /* synthesis syn_keep=1 */ ;
wire out144 /* synthesis syn_keep=1 */ ;
wire out145 /* synthesis syn_keep=1 */ ;
wire out146 /* synthesis syn_keep=1 */ ;
wire out147 /* synthesis syn_keep=1 */ ;
wire out148 /* synthesis syn_keep=1 */ ;
wire out149 /* synthesis syn_keep=1 */ ;
wire out150 /* synthesis syn_keep=1 */ ;
wire out151 /* synthesis syn_keep=1 */ ;
wire out152 /* synthesis syn_keep=1 */ ;
wire out153 /* synthesis syn_keep=1 */ ;
wire out154 /* synthesis syn_keep=1 */ ;
wire out155 /* synthesis syn_keep=1 */ ;
wire out156 /* synthesis syn_keep=1 */ ;
wire out157 /* synthesis syn_keep=1 */ ;
wire out158 /* synthesis syn_keep=1 */ ;
wire out159 /* synthesis syn_keep=1 */ ;
wire out160 /* synthesis syn_keep=1 */ ;
wire out161 /* synthesis syn_keep=1 */ ;
wire out162 /* synthesis syn_keep=1 */ ;
wire out163 /* synthesis syn_keep=1 */ ;
wire out164 /* synthesis syn_keep=1 */ ;
wire out165 /* synthesis syn_keep=1 */ ;
wire out166 /* synthesis syn_keep=1 */ ;
wire out167 /* synthesis syn_keep=1 */ ;
wire out168 /* synthesis syn_keep=1 */ ;
wire out169 /* synthesis syn_keep=1 */ ;
wire out170 /* synthesis syn_keep=1 */ ;
wire out171 /* synthesis syn_keep=1 */ ;
wire out172 /* synthesis syn_keep=1 */ ;
wire out173 /* synthesis syn_keep=1 */ ;
wire out174 /* synthesis syn_keep=1 */ ;
wire out175 /* synthesis syn_keep=1 */ ;
wire out176 /* synthesis syn_keep=1 */ ;
wire out177 /* synthesis syn_keep=1 */ ;
wire out178 /* synthesis syn_keep=1 */ ;
wire out179 /* synthesis syn_keep=1 */ ;
wire out180 /* synthesis syn_keep=1 */ ;
wire out181 /* synthesis syn_keep=1 */ ;
wire out182 /* synthesis syn_keep=1 */ ;
wire out183 /* synthesis syn_keep=1 */ ;
wire out184 /* synthesis syn_keep=1 */ ;
wire out185 /* synthesis syn_keep=1 */ ;
wire out186 /* synthesis syn_keep=1 */ ;
wire out187 /* synthesis syn_keep=1 */ ;
wire out188 /* synthesis syn_keep=1 */ ;
wire out189 /* synthesis syn_keep=1 */ ;
wire out190 /* synthesis syn_keep=1 */ ;
wire out191 /* synthesis syn_keep=1 */ ;
wire out192 /* synthesis syn_keep=1 */ ;
wire out193 /* synthesis syn_keep=1 */ ;
wire out194 /* synthesis syn_keep=1 */ ;
wire out195 /* synthesis syn_keep=1 */ ;
wire out196 /* synthesis syn_keep=1 */ ;
wire out197 /* synthesis syn_keep=1 */ ;
wire out198 /* synthesis syn_keep=1 */ ;
wire out199 /* synthesis syn_keep=1 */ ;
wire out200 /* synthesis syn_keep=1 */ ;
wire out201 /* synthesis syn_keep=1 */ ;
wire out202 /* synthesis syn_keep=1 */ ;
wire out203 /* synthesis syn_keep=1 */ ;
wire out204 /* synthesis syn_keep=1 */ ;
wire out205 /* synthesis syn_keep=1 */ ;
wire out206 /* synthesis syn_keep=1 */ ;
wire out207 /* synthesis syn_keep=1 */ ;
wire out208 /* synthesis syn_keep=1 */ ;
wire out209 /* synthesis syn_keep=1 */ ;
wire out210 /* synthesis syn_keep=1 */ ;
wire out211 /* synthesis syn_keep=1 */ ;
wire out212 /* synthesis syn_keep=1 */ ;
wire out213 /* synthesis syn_keep=1 */ ;
wire out214 /* synthesis syn_keep=1 */ ;
wire out215 /* synthesis syn_keep=1 */ ;
wire out216 /* synthesis syn_keep=1 */ ;
wire out217 /* synthesis syn_keep=1 */ ;
wire out218 /* synthesis syn_keep=1 */ ;
wire out219 /* synthesis syn_keep=1 */ ;
wire out220 /* synthesis syn_keep=1 */ ;
wire out221 /* synthesis syn_keep=1 */ ;
wire out222 /* synthesis syn_keep=1 */ ;
wire out223 /* synthesis syn_keep=1 */ ;
wire out224 /* synthesis syn_keep=1 */ ;
wire out225 /* synthesis syn_keep=1 */ ;
wire out226 /* synthesis syn_keep=1 */ ;
wire out227 /* synthesis syn_keep=1 */ ;
wire out228 /* synthesis syn_keep=1 */ ;
wire out229 /* synthesis syn_keep=1 */ ;
wire out230 /* synthesis syn_keep=1 */ ;
wire out231 /* synthesis syn_keep=1 */ ;
wire out232 /* synthesis syn_keep=1 */ ;
wire out233 /* synthesis syn_keep=1 */ ;
wire out234 /* synthesis syn_keep=1 */ ;
wire out235 /* synthesis syn_keep=1 */ ;
wire out236 /* synthesis syn_keep=1 */ ;
wire out237 /* synthesis syn_keep=1 */ ;
wire out238 /* synthesis syn_keep=1 */ ;
wire out239 /* synthesis syn_keep=1 */ ;
wire out240 /* synthesis syn_keep=1 */ ;
wire out241 /* synthesis syn_keep=1 */ ;
wire out242 /* synthesis syn_keep=1 */ ;
wire out243 /* synthesis syn_keep=1 */ ;
wire out244 /* synthesis syn_keep=1 */ ;
wire out245 /* synthesis syn_keep=1 */ ;
wire out246 /* synthesis syn_keep=1 */ ;
wire out247 /* synthesis syn_keep=1 */ ;
wire out248 /* synthesis syn_keep=1 */ ;
wire out249 /* synthesis syn_keep=1 */ ;
wire out250 /* synthesis syn_keep=1 */ ;
wire out251 /* synthesis syn_keep=1 */ ;
wire out252 /* synthesis syn_keep=1 */ ;
wire out253 /* synthesis syn_keep=1 */ ;
wire out254 /* synthesis syn_keep=1 */ ;

del_elem_v2 inst0(
.clk(clk),
.delay_in(start),
.delay_out(out0),
.reg_out(regs_out[0])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst1(
.clk(clk),
.delay_in(out0),
.delay_out(out1),
.reg_out(regs_out[1])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst2(
.clk(clk),
.delay_in(out1),
.delay_out(out2),
.reg_out(regs_out[2])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst3(
.clk(clk),
.delay_in(out2),
.delay_out(out3),
.reg_out(regs_out[3])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst4(
.clk(clk),
.delay_in(out3),
.delay_out(out4),
.reg_out(regs_out[4])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst5(
.clk(clk),
.delay_in(out4),
.delay_out(out5),
.reg_out(regs_out[5])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst6(
.clk(clk),
.delay_in(out5),
.delay_out(out6),
.reg_out(regs_out[6])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst7(
.clk(clk),
.delay_in(out6),
.delay_out(out7),
.reg_out(regs_out[7])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst8(
.clk(clk),
.delay_in(out7),
.delay_out(out8),
.reg_out(regs_out[8])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst9(
.clk(clk),
.delay_in(out8),
.delay_out(out9),
.reg_out(regs_out[9])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst10(
.clk(clk),
.delay_in(out9),
.delay_out(out10),
.reg_out(regs_out[10])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst11(
.clk(clk),
.delay_in(out10),
.delay_out(out11),
.reg_out(regs_out[11])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst12(
.clk(clk),
.delay_in(out11),
.delay_out(out12),
.reg_out(regs_out[12])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst13(
.clk(clk),
.delay_in(out12),
.delay_out(out13),
.reg_out(regs_out[13])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst14(
.clk(clk),
.delay_in(out13),
.delay_out(out14),
.reg_out(regs_out[14])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst15(
.clk(clk),
.delay_in(out14),
.delay_out(out15),
.reg_out(regs_out[15])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst16(
.clk(clk),
.delay_in(out15),
.delay_out(out16),
.reg_out(regs_out[16])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst17(
.clk(clk),
.delay_in(out16),
.delay_out(out17),
.reg_out(regs_out[17])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst18(
.clk(clk),
.delay_in(out17),
.delay_out(out18),
.reg_out(regs_out[18])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst19(
.clk(clk),
.delay_in(out18),
.delay_out(out19),
.reg_out(regs_out[19])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst20(
.clk(clk),
.delay_in(out19),
.delay_out(out20),
.reg_out(regs_out[20])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst21(
.clk(clk),
.delay_in(out20),
.delay_out(out21),
.reg_out(regs_out[21])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst22(
.clk(clk),
.delay_in(out21),
.delay_out(out22),
.reg_out(regs_out[22])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst23(
.clk(clk),
.delay_in(out22),
.delay_out(out23),
.reg_out(regs_out[23])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst24(
.clk(clk),
.delay_in(out23),
.delay_out(out24),
.reg_out(regs_out[24])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst25(
.clk(clk),
.delay_in(out24),
.delay_out(out25),
.reg_out(regs_out[25])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst26(
.clk(clk),
.delay_in(out25),
.delay_out(out26),
.reg_out(regs_out[26])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst27(
.clk(clk),
.delay_in(out26),
.delay_out(out27),
.reg_out(regs_out[27])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst28(
.clk(clk),
.delay_in(out27),
.delay_out(out28),
.reg_out(regs_out[28])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst29(
.clk(clk),
.delay_in(out28),
.delay_out(out29),
.reg_out(regs_out[29])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst30(
.clk(clk),
.delay_in(out29),
.delay_out(out30),
.reg_out(regs_out[30])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst31(
.clk(clk),
.delay_in(out30),
.delay_out(out31),
.reg_out(regs_out[31])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst32(
.clk(clk),
.delay_in(out31),
.delay_out(out32),
.reg_out(regs_out[32])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst33(
.clk(clk),
.delay_in(out32),
.delay_out(out33),
.reg_out(regs_out[33])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst34(
.clk(clk),
.delay_in(out33),
.delay_out(out34),
.reg_out(regs_out[34])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst35(
.clk(clk),
.delay_in(out34),
.delay_out(out35),
.reg_out(regs_out[35])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst36(
.clk(clk),
.delay_in(out35),
.delay_out(out36),
.reg_out(regs_out[36])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst37(
.clk(clk),
.delay_in(out36),
.delay_out(out37),
.reg_out(regs_out[37])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst38(
.clk(clk),
.delay_in(out37),
.delay_out(out38),
.reg_out(regs_out[38])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst39(
.clk(clk),
.delay_in(out38),
.delay_out(out39),
.reg_out(regs_out[39])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst40(
.clk(clk),
.delay_in(out39),
.delay_out(out40),
.reg_out(regs_out[40])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst41(
.clk(clk),
.delay_in(out40),
.delay_out(out41),
.reg_out(regs_out[41])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst42(
.clk(clk),
.delay_in(out41),
.delay_out(out42),
.reg_out(regs_out[42])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst43(
.clk(clk),
.delay_in(out42),
.delay_out(out43),
.reg_out(regs_out[43])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst44(
.clk(clk),
.delay_in(out43),
.delay_out(out44),
.reg_out(regs_out[44])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst45(
.clk(clk),
.delay_in(out44),
.delay_out(out45),
.reg_out(regs_out[45])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst46(
.clk(clk),
.delay_in(out45),
.delay_out(out46),
.reg_out(regs_out[46])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst47(
.clk(clk),
.delay_in(out46),
.delay_out(out47),
.reg_out(regs_out[47])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst48(
.clk(clk),
.delay_in(out47),
.delay_out(out48),
.reg_out(regs_out[48])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst49(
.clk(clk),
.delay_in(out48),
.delay_out(out49),
.reg_out(regs_out[49])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst50(
.clk(clk),
.delay_in(out49),
.delay_out(out50),
.reg_out(regs_out[50])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst51(
.clk(clk),
.delay_in(out50),
.delay_out(out51),
.reg_out(regs_out[51])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst52(
.clk(clk),
.delay_in(out51),
.delay_out(out52),
.reg_out(regs_out[52])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst53(
.clk(clk),
.delay_in(out52),
.delay_out(out53),
.reg_out(regs_out[53])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst54(
.clk(clk),
.delay_in(out53),
.delay_out(out54),
.reg_out(regs_out[54])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst55(
.clk(clk),
.delay_in(out54),
.delay_out(out55),
.reg_out(regs_out[55])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst56(
.clk(clk),
.delay_in(out55),
.delay_out(out56),
.reg_out(regs_out[56])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst57(
.clk(clk),
.delay_in(out56),
.delay_out(out57),
.reg_out(regs_out[57])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst58(
.clk(clk),
.delay_in(out57),
.delay_out(out58),
.reg_out(regs_out[58])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst59(
.clk(clk),
.delay_in(out58),
.delay_out(out59),
.reg_out(regs_out[59])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst60(
.clk(clk),
.delay_in(out59),
.delay_out(out60),
.reg_out(regs_out[60])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst61(
.clk(clk),
.delay_in(out60),
.delay_out(out61),
.reg_out(regs_out[61])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst62(
.clk(clk),
.delay_in(out61),
.delay_out(out62),
.reg_out(regs_out[62])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst63(
.clk(clk),
.delay_in(out62),
.delay_out(out63),
.reg_out(regs_out[63])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst64(
.clk(clk),
.delay_in(out63),
.delay_out(out64),
.reg_out(regs_out[64])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst65(
.clk(clk),
.delay_in(out64),
.delay_out(out65),
.reg_out(regs_out[65])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst66(
.clk(clk),
.delay_in(out65),
.delay_out(out66),
.reg_out(regs_out[66])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst67(
.clk(clk),
.delay_in(out66),
.delay_out(out67),
.reg_out(regs_out[67])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst68(
.clk(clk),
.delay_in(out67),
.delay_out(out68),
.reg_out(regs_out[68])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst69(
.clk(clk),
.delay_in(out68),
.delay_out(out69),
.reg_out(regs_out[69])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst70(
.clk(clk),
.delay_in(out69),
.delay_out(out70),
.reg_out(regs_out[70])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst71(
.clk(clk),
.delay_in(out70),
.delay_out(out71),
.reg_out(regs_out[71])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst72(
.clk(clk),
.delay_in(out71),
.delay_out(out72),
.reg_out(regs_out[72])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst73(
.clk(clk),
.delay_in(out72),
.delay_out(out73),
.reg_out(regs_out[73])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst74(
.clk(clk),
.delay_in(out73),
.delay_out(out74),
.reg_out(regs_out[74])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst75(
.clk(clk),
.delay_in(out74),
.delay_out(out75),
.reg_out(regs_out[75])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst76(
.clk(clk),
.delay_in(out75),
.delay_out(out76),
.reg_out(regs_out[76])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst77(
.clk(clk),
.delay_in(out76),
.delay_out(out77),
.reg_out(regs_out[77])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst78(
.clk(clk),
.delay_in(out77),
.delay_out(out78),
.reg_out(regs_out[78])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst79(
.clk(clk),
.delay_in(out78),
.delay_out(out79),
.reg_out(regs_out[79])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst80(
.clk(clk),
.delay_in(out79),
.delay_out(out80),
.reg_out(regs_out[80])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst81(
.clk(clk),
.delay_in(out80),
.delay_out(out81),
.reg_out(regs_out[81])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst82(
.clk(clk),
.delay_in(out81),
.delay_out(out82),
.reg_out(regs_out[82])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst83(
.clk(clk),
.delay_in(out82),
.delay_out(out83),
.reg_out(regs_out[83])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst84(
.clk(clk),
.delay_in(out83),
.delay_out(out84),
.reg_out(regs_out[84])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst85(
.clk(clk),
.delay_in(out84),
.delay_out(out85),
.reg_out(regs_out[85])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst86(
.clk(clk),
.delay_in(out85),
.delay_out(out86),
.reg_out(regs_out[86])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst87(
.clk(clk),
.delay_in(out86),
.delay_out(out87),
.reg_out(regs_out[87])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst88(
.clk(clk),
.delay_in(out87),
.delay_out(out88),
.reg_out(regs_out[88])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst89(
.clk(clk),
.delay_in(out88),
.delay_out(out89),
.reg_out(regs_out[89])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst90(
.clk(clk),
.delay_in(out89),
.delay_out(out90),
.reg_out(regs_out[90])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst91(
.clk(clk),
.delay_in(out90),
.delay_out(out91),
.reg_out(regs_out[91])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst92(
.clk(clk),
.delay_in(out91),
.delay_out(out92),
.reg_out(regs_out[92])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst93(
.clk(clk),
.delay_in(out92),
.delay_out(out93),
.reg_out(regs_out[93])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst94(
.clk(clk),
.delay_in(out93),
.delay_out(out94),
.reg_out(regs_out[94])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst95(
.clk(clk),
.delay_in(out94),
.delay_out(out95),
.reg_out(regs_out[95])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst96(
.clk(clk),
.delay_in(out95),
.delay_out(out96),
.reg_out(regs_out[96])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst97(
.clk(clk),
.delay_in(out96),
.delay_out(out97),
.reg_out(regs_out[97])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst98(
.clk(clk),
.delay_in(out97),
.delay_out(out98),
.reg_out(regs_out[98])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst99(
.clk(clk),
.delay_in(out98),
.delay_out(out99),
.reg_out(regs_out[99])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst100(
.clk(clk),
.delay_in(out99),
.delay_out(out100),
.reg_out(regs_out[100])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst101(
.clk(clk),
.delay_in(out100),
.delay_out(out101),
.reg_out(regs_out[101])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst102(
.clk(clk),
.delay_in(out101),
.delay_out(out102),
.reg_out(regs_out[102])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst103(
.clk(clk),
.delay_in(out102),
.delay_out(out103),
.reg_out(regs_out[103])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst104(
.clk(clk),
.delay_in(out103),
.delay_out(out104),
.reg_out(regs_out[104])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst105(
.clk(clk),
.delay_in(out104),
.delay_out(out105),
.reg_out(regs_out[105])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst106(
.clk(clk),
.delay_in(out105),
.delay_out(out106),
.reg_out(regs_out[106])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst107(
.clk(clk),
.delay_in(out106),
.delay_out(out107),
.reg_out(regs_out[107])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst108(
.clk(clk),
.delay_in(out107),
.delay_out(out108),
.reg_out(regs_out[108])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst109(
.clk(clk),
.delay_in(out108),
.delay_out(out109),
.reg_out(regs_out[109])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst110(
.clk(clk),
.delay_in(out109),
.delay_out(out110),
.reg_out(regs_out[110])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst111(
.clk(clk),
.delay_in(out110),
.delay_out(out111),
.reg_out(regs_out[111])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst112(
.clk(clk),
.delay_in(out111),
.delay_out(out112),
.reg_out(regs_out[112])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst113(
.clk(clk),
.delay_in(out112),
.delay_out(out113),
.reg_out(regs_out[113])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst114(
.clk(clk),
.delay_in(out113),
.delay_out(out114),
.reg_out(regs_out[114])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst115(
.clk(clk),
.delay_in(out114),
.delay_out(out115),
.reg_out(regs_out[115])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst116(
.clk(clk),
.delay_in(out115),
.delay_out(out116),
.reg_out(regs_out[116])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst117(
.clk(clk),
.delay_in(out116),
.delay_out(out117),
.reg_out(regs_out[117])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst118(
.clk(clk),
.delay_in(out117),
.delay_out(out118),
.reg_out(regs_out[118])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst119(
.clk(clk),
.delay_in(out118),
.delay_out(out119),
.reg_out(regs_out[119])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst120(
.clk(clk),
.delay_in(out119),
.delay_out(out120),
.reg_out(regs_out[120])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst121(
.clk(clk),
.delay_in(out120),
.delay_out(out121),
.reg_out(regs_out[121])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst122(
.clk(clk),
.delay_in(out121),
.delay_out(out122),
.reg_out(regs_out[122])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst123(
.clk(clk),
.delay_in(out122),
.delay_out(out123),
.reg_out(regs_out[123])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst124(
.clk(clk),
.delay_in(out123),
.delay_out(out124),
.reg_out(regs_out[124])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst125(
.clk(clk),
.delay_in(out124),
.delay_out(out125),
.reg_out(regs_out[125])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst126(
.clk(clk),
.delay_in(out125),
.delay_out(out126),
.reg_out(regs_out[126])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst127(
.clk(clk),
.delay_in(out126),
.delay_out(out127),
.reg_out(regs_out[127])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst128(
.clk(clk),
.delay_in(out127),
.delay_out(out128),
.reg_out(regs_out[128])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst129(
.clk(clk),
.delay_in(out128),
.delay_out(out129),
.reg_out(regs_out[129])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst130(
.clk(clk),
.delay_in(out129),
.delay_out(out130),
.reg_out(regs_out[130])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst131(
.clk(clk),
.delay_in(out130),
.delay_out(out131),
.reg_out(regs_out[131])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst132(
.clk(clk),
.delay_in(out131),
.delay_out(out132),
.reg_out(regs_out[132])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst133(
.clk(clk),
.delay_in(out132),
.delay_out(out133),
.reg_out(regs_out[133])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst134(
.clk(clk),
.delay_in(out133),
.delay_out(out134),
.reg_out(regs_out[134])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst135(
.clk(clk),
.delay_in(out134),
.delay_out(out135),
.reg_out(regs_out[135])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst136(
.clk(clk),
.delay_in(out135),
.delay_out(out136),
.reg_out(regs_out[136])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst137(
.clk(clk),
.delay_in(out136),
.delay_out(out137),
.reg_out(regs_out[137])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst138(
.clk(clk),
.delay_in(out137),
.delay_out(out138),
.reg_out(regs_out[138])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst139(
.clk(clk),
.delay_in(out138),
.delay_out(out139),
.reg_out(regs_out[139])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst140(
.clk(clk),
.delay_in(out139),
.delay_out(out140),
.reg_out(regs_out[140])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst141(
.clk(clk),
.delay_in(out140),
.delay_out(out141),
.reg_out(regs_out[141])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst142(
.clk(clk),
.delay_in(out141),
.delay_out(out142),
.reg_out(regs_out[142])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst143(
.clk(clk),
.delay_in(out142),
.delay_out(out143),
.reg_out(regs_out[143])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst144(
.clk(clk),
.delay_in(out143),
.delay_out(out144),
.reg_out(regs_out[144])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst145(
.clk(clk),
.delay_in(out144),
.delay_out(out145),
.reg_out(regs_out[145])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst146(
.clk(clk),
.delay_in(out145),
.delay_out(out146),
.reg_out(regs_out[146])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst147(
.clk(clk),
.delay_in(out146),
.delay_out(out147),
.reg_out(regs_out[147])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst148(
.clk(clk),
.delay_in(out147),
.delay_out(out148),
.reg_out(regs_out[148])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst149(
.clk(clk),
.delay_in(out148),
.delay_out(out149),
.reg_out(regs_out[149])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst150(
.clk(clk),
.delay_in(out149),
.delay_out(out150),
.reg_out(regs_out[150])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst151(
.clk(clk),
.delay_in(out150),
.delay_out(out151),
.reg_out(regs_out[151])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst152(
.clk(clk),
.delay_in(out151),
.delay_out(out152),
.reg_out(regs_out[152])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst153(
.clk(clk),
.delay_in(out152),
.delay_out(out153),
.reg_out(regs_out[153])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst154(
.clk(clk),
.delay_in(out153),
.delay_out(out154),
.reg_out(regs_out[154])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst155(
.clk(clk),
.delay_in(out154),
.delay_out(out155),
.reg_out(regs_out[155])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst156(
.clk(clk),
.delay_in(out155),
.delay_out(out156),
.reg_out(regs_out[156])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst157(
.clk(clk),
.delay_in(out156),
.delay_out(out157),
.reg_out(regs_out[157])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst158(
.clk(clk),
.delay_in(out157),
.delay_out(out158),
.reg_out(regs_out[158])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst159(
.clk(clk),
.delay_in(out158),
.delay_out(out159),
.reg_out(regs_out[159])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst160(
.clk(clk),
.delay_in(out159),
.delay_out(out160),
.reg_out(regs_out[160])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst161(
.clk(clk),
.delay_in(out160),
.delay_out(out161),
.reg_out(regs_out[161])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst162(
.clk(clk),
.delay_in(out161),
.delay_out(out162),
.reg_out(regs_out[162])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst163(
.clk(clk),
.delay_in(out162),
.delay_out(out163),
.reg_out(regs_out[163])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst164(
.clk(clk),
.delay_in(out163),
.delay_out(out164),
.reg_out(regs_out[164])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst165(
.clk(clk),
.delay_in(out164),
.delay_out(out165),
.reg_out(regs_out[165])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst166(
.clk(clk),
.delay_in(out165),
.delay_out(out166),
.reg_out(regs_out[166])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst167(
.clk(clk),
.delay_in(out166),
.delay_out(out167),
.reg_out(regs_out[167])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst168(
.clk(clk),
.delay_in(out167),
.delay_out(out168),
.reg_out(regs_out[168])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst169(
.clk(clk),
.delay_in(out168),
.delay_out(out169),
.reg_out(regs_out[169])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst170(
.clk(clk),
.delay_in(out169),
.delay_out(out170),
.reg_out(regs_out[170])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst171(
.clk(clk),
.delay_in(out170),
.delay_out(out171),
.reg_out(regs_out[171])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst172(
.clk(clk),
.delay_in(out171),
.delay_out(out172),
.reg_out(regs_out[172])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst173(
.clk(clk),
.delay_in(out172),
.delay_out(out173),
.reg_out(regs_out[173])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst174(
.clk(clk),
.delay_in(out173),
.delay_out(out174),
.reg_out(regs_out[174])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst175(
.clk(clk),
.delay_in(out174),
.delay_out(out175),
.reg_out(regs_out[175])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst176(
.clk(clk),
.delay_in(out175),
.delay_out(out176),
.reg_out(regs_out[176])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst177(
.clk(clk),
.delay_in(out176),
.delay_out(out177),
.reg_out(regs_out[177])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst178(
.clk(clk),
.delay_in(out177),
.delay_out(out178),
.reg_out(regs_out[178])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst179(
.clk(clk),
.delay_in(out178),
.delay_out(out179),
.reg_out(regs_out[179])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst180(
.clk(clk),
.delay_in(out179),
.delay_out(out180),
.reg_out(regs_out[180])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst181(
.clk(clk),
.delay_in(out180),
.delay_out(out181),
.reg_out(regs_out[181])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst182(
.clk(clk),
.delay_in(out181),
.delay_out(out182),
.reg_out(regs_out[182])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst183(
.clk(clk),
.delay_in(out182),
.delay_out(out183),
.reg_out(regs_out[183])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst184(
.clk(clk),
.delay_in(out183),
.delay_out(out184),
.reg_out(regs_out[184])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst185(
.clk(clk),
.delay_in(out184),
.delay_out(out185),
.reg_out(regs_out[185])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst186(
.clk(clk),
.delay_in(out185),
.delay_out(out186),
.reg_out(regs_out[186])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst187(
.clk(clk),
.delay_in(out186),
.delay_out(out187),
.reg_out(regs_out[187])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst188(
.clk(clk),
.delay_in(out187),
.delay_out(out188),
.reg_out(regs_out[188])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst189(
.clk(clk),
.delay_in(out188),
.delay_out(out189),
.reg_out(regs_out[189])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst190(
.clk(clk),
.delay_in(out189),
.delay_out(out190),
.reg_out(regs_out[190])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst191(
.clk(clk),
.delay_in(out190),
.delay_out(out191),
.reg_out(regs_out[191])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst192(
.clk(clk),
.delay_in(out191),
.delay_out(out192),
.reg_out(regs_out[192])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst193(
.clk(clk),
.delay_in(out192),
.delay_out(out193),
.reg_out(regs_out[193])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst194(
.clk(clk),
.delay_in(out193),
.delay_out(out194),
.reg_out(regs_out[194])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst195(
.clk(clk),
.delay_in(out194),
.delay_out(out195),
.reg_out(regs_out[195])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst196(
.clk(clk),
.delay_in(out195),
.delay_out(out196),
.reg_out(regs_out[196])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst197(
.clk(clk),
.delay_in(out196),
.delay_out(out197),
.reg_out(regs_out[197])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst198(
.clk(clk),
.delay_in(out197),
.delay_out(out198),
.reg_out(regs_out[198])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst199(
.clk(clk),
.delay_in(out198),
.delay_out(out199),
.reg_out(regs_out[199])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst200(
.clk(clk),
.delay_in(out199),
.delay_out(out200),
.reg_out(regs_out[200])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst201(
.clk(clk),
.delay_in(out200),
.delay_out(out201),
.reg_out(regs_out[201])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst202(
.clk(clk),
.delay_in(out201),
.delay_out(out202),
.reg_out(regs_out[202])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst203(
.clk(clk),
.delay_in(out202),
.delay_out(out203),
.reg_out(regs_out[203])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst204(
.clk(clk),
.delay_in(out203),
.delay_out(out204),
.reg_out(regs_out[204])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst205(
.clk(clk),
.delay_in(out204),
.delay_out(out205),
.reg_out(regs_out[205])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst206(
.clk(clk),
.delay_in(out205),
.delay_out(out206),
.reg_out(regs_out[206])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst207(
.clk(clk),
.delay_in(out206),
.delay_out(out207),
.reg_out(regs_out[207])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst208(
.clk(clk),
.delay_in(out207),
.delay_out(out208),
.reg_out(regs_out[208])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst209(
.clk(clk),
.delay_in(out208),
.delay_out(out209),
.reg_out(regs_out[209])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst210(
.clk(clk),
.delay_in(out209),
.delay_out(out210),
.reg_out(regs_out[210])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst211(
.clk(clk),
.delay_in(out210),
.delay_out(out211),
.reg_out(regs_out[211])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst212(
.clk(clk),
.delay_in(out211),
.delay_out(out212),
.reg_out(regs_out[212])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst213(
.clk(clk),
.delay_in(out212),
.delay_out(out213),
.reg_out(regs_out[213])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst214(
.clk(clk),
.delay_in(out213),
.delay_out(out214),
.reg_out(regs_out[214])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst215(
.clk(clk),
.delay_in(out214),
.delay_out(out215),
.reg_out(regs_out[215])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst216(
.clk(clk),
.delay_in(out215),
.delay_out(out216),
.reg_out(regs_out[216])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst217(
.clk(clk),
.delay_in(out216),
.delay_out(out217),
.reg_out(regs_out[217])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst218(
.clk(clk),
.delay_in(out217),
.delay_out(out218),
.reg_out(regs_out[218])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst219(
.clk(clk),
.delay_in(out218),
.delay_out(out219),
.reg_out(regs_out[219])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst220(
.clk(clk),
.delay_in(out219),
.delay_out(out220),
.reg_out(regs_out[220])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst221(
.clk(clk),
.delay_in(out220),
.delay_out(out221),
.reg_out(regs_out[221])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst222(
.clk(clk),
.delay_in(out221),
.delay_out(out222),
.reg_out(regs_out[222])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst223(
.clk(clk),
.delay_in(out222),
.delay_out(out223),
.reg_out(regs_out[223])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst224(
.clk(clk),
.delay_in(out223),
.delay_out(out224),
.reg_out(regs_out[224])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst225(
.clk(clk),
.delay_in(out224),
.delay_out(out225),
.reg_out(regs_out[225])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst226(
.clk(clk),
.delay_in(out225),
.delay_out(out226),
.reg_out(regs_out[226])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst227(
.clk(clk),
.delay_in(out226),
.delay_out(out227),
.reg_out(regs_out[227])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst228(
.clk(clk),
.delay_in(out227),
.delay_out(out228),
.reg_out(regs_out[228])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst229(
.clk(clk),
.delay_in(out228),
.delay_out(out229),
.reg_out(regs_out[229])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst230(
.clk(clk),
.delay_in(out229),
.delay_out(out230),
.reg_out(regs_out[230])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst231(
.clk(clk),
.delay_in(out230),
.delay_out(out231),
.reg_out(regs_out[231])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst232(
.clk(clk),
.delay_in(out231),
.delay_out(out232),
.reg_out(regs_out[232])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst233(
.clk(clk),
.delay_in(out232),
.delay_out(out233),
.reg_out(regs_out[233])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst234(
.clk(clk),
.delay_in(out233),
.delay_out(out234),
.reg_out(regs_out[234])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst235(
.clk(clk),
.delay_in(out234),
.delay_out(out235),
.reg_out(regs_out[235])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst236(
.clk(clk),
.delay_in(out235),
.delay_out(out236),
.reg_out(regs_out[236])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst237(
.clk(clk),
.delay_in(out236),
.delay_out(out237),
.reg_out(regs_out[237])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst238(
.clk(clk),
.delay_in(out237),
.delay_out(out238),
.reg_out(regs_out[238])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst239(
.clk(clk),
.delay_in(out238),
.delay_out(out239),
.reg_out(regs_out[239])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst240(
.clk(clk),
.delay_in(out239),
.delay_out(out240),
.reg_out(regs_out[240])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst241(
.clk(clk),
.delay_in(out240),
.delay_out(out241),
.reg_out(regs_out[241])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst242(
.clk(clk),
.delay_in(out241),
.delay_out(out242),
.reg_out(regs_out[242])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst243(
.clk(clk),
.delay_in(out242),
.delay_out(out243),
.reg_out(regs_out[243])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst244(
.clk(clk),
.delay_in(out243),
.delay_out(out244),
.reg_out(regs_out[244])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst245(
.clk(clk),
.delay_in(out244),
.delay_out(out245),
.reg_out(regs_out[245])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst246(
.clk(clk),
.delay_in(out245),
.delay_out(out246),
.reg_out(regs_out[246])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst247(
.clk(clk),
.delay_in(out246),
.delay_out(out247),
.reg_out(regs_out[247])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst248(
.clk(clk),
.delay_in(out247),
.delay_out(out248),
.reg_out(regs_out[248])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst249(
.clk(clk),
.delay_in(out248),
.delay_out(out249),
.reg_out(regs_out[249])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst250(
.clk(clk),
.delay_in(out249),
.delay_out(out250),
.reg_out(regs_out[250])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst251(
.clk(clk),
.delay_in(out250),
.delay_out(out251),
.reg_out(regs_out[251])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst252(
.clk(clk),
.delay_in(out251),
.delay_out(out252),
.reg_out(regs_out[252])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst253(
.clk(clk),
.delay_in(out252),
.delay_out(out253),
.reg_out(regs_out[253])
) /* synthesis syn_noprune=1 */;

del_elem_v2 inst254(
.clk(clk),
.delay_in(out253),
.delay_out(out254),
.reg_out(regs_out[254])
) /* synthesis syn_noprune=1 */;

assign out = out254;

endmodule
